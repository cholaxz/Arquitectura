`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:38:03 10/08/2018 
// Design Name: 
// Module Name:    program_memory 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module program_memory#(
	parameter ADDR_LENGTH = 11,
	parameter DATA_LENGTH = 16,
	parameter program = "/home/agustin/Desktop/Arquitectura/TP3/code/program.bin"
)(
	input clk,
	input [ADDR_LENGTH - 1 : 0]addr,
	input Wr,
	input[DATA_LENGTH - 1 : 0] inData,
	output reg[DATA_LENGTH - 1 : 0] instruction
   );
	
	localparam MEM_SIZE = 2 ^ ADDR_LENGTH ;
	reg [DATA_LENGTH - 1 : 0]memory[0 : MEM_SIZE];
	
	
	initial begin
	if(program != "")
		$readmemb(program, memory);
	else
		begin
			memory[0] = 16'b0001000000000001; //Load Addr1
			memory[1] = 16'b0010000000000010; //Add Acc + Addr2
			memory[2] = 16'b0000100000000000; //Store Acc in Addr0
			memory[3] = 16'b0000000000000000; //Halt
		end
	end

always @(posedge clk)
begin
	if(Wr == 1)
		memory[addr] <= inData;
	else
		instruction <= memory[addr];
end



endmodule